library verilog;
use verilog.vl_types.all;
entity temporizador_vlg_vec_tst is
end temporizador_vlg_vec_tst;
