library verilog;
use verilog.vl_types.all;
entity Luces_vlg_vec_tst is
end Luces_vlg_vec_tst;
