library verilog;
use verilog.vl_types.all;
entity minutos_vlg_vec_tst is
end minutos_vlg_vec_tst;
