library verilog;
use verilog.vl_types.all;
entity contador_3_vlg_check_tst is
    port(
        ADES            : in     vl_logic;
        ADM             : in     vl_logic;
        ADS             : in     vl_logic;
        AUM             : in     vl_logic;
        AUS             : in     vl_logic;
        BDES            : in     vl_logic;
        BDM             : in     vl_logic;
        BDS             : in     vl_logic;
        BUM             : in     vl_logic;
        \BUS\           : in     vl_logic;
        CDES            : in     vl_logic;
        CDM             : in     vl_logic;
        CDS             : in     vl_logic;
        CUM             : in     vl_logic;
        CUS             : in     vl_logic;
        DDES            : in     vl_logic;
        DDM             : in     vl_logic;
        DDS             : in     vl_logic;
        DUM             : in     vl_logic;
        DUS             : in     vl_logic;
        EDES            : in     vl_logic;
        EDM             : in     vl_logic;
        EDS             : in     vl_logic;
        EUM             : in     vl_logic;
        EUS             : in     vl_logic;
        FDES            : in     vl_logic;
        FDM             : in     vl_logic;
        FDS             : in     vl_logic;
        FUM             : in     vl_logic;
        FUS             : in     vl_logic;
        GDES            : in     vl_logic;
        GDM             : in     vl_logic;
        GDS             : in     vl_logic;
        GUM             : in     vl_logic;
        GUS             : in     vl_logic;
        \OUT\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end contador_3_vlg_check_tst;
