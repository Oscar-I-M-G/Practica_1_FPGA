library verilog;
use verilog.vl_types.all;
entity temporizador_50MHz_vlg_vec_tst is
end temporizador_50MHz_vlg_vec_tst;
