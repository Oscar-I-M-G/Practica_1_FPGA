library verilog;
use verilog.vl_types.all;
entity Conversor_vlg_vec_tst is
end Conversor_vlg_vec_tst;
