library verilog;
use verilog.vl_types.all;
entity contador_2_vlg_vec_tst is
end contador_2_vlg_vec_tst;
