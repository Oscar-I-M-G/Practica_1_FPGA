library verilog;
use verilog.vl_types.all;
entity temporizador_50MHz_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end temporizador_50MHz_vlg_check_tst;
